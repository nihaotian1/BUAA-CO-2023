`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:40:55 11/09/2023 
// Design Name: 
// Module Name:    W 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module W(
    input clk,
    input reset,
    input [31:0] Instr_M,
    input [31:0] pc_M,
    input [31:0] pc4_M,
    input [31:0] outC_M,
    input [31:0] ReadData_M,
    input [3:0] Tnew_M,
    output [31:0] Instr_W,
    output [31:0] pc_W,
    output [31:0] pc4_W,
    output [31:0] ReadData_W,
    output [31:0] outC_W,
    output [3:0] Tnew_W
    );

    reg [31:0] Instr;
    reg [31:0] pc;
    reg [31:0] pc4;
    reg [31:0] outC;
    reg [31:0] ReadData;
    reg [3:0] Tnew;

    always @(posedge clk) begin
        if(reset == 1'b1) begin
            Instr <= 32'h0000_0000;
            pc <= 32'h0000_0000;
            pc4 <= 32'h0000_0000;
            outC <= 32'h0000_0000;
            ReadData <= 32'h0000_0000;
            Tnew <= 4'h0;
        end
        else begin
            Instr <= Instr_M;
            pc <= pc_M;
            pc4 <= pc4_M;
            outC <= outC_M;
            ReadData <= ReadData_M;
            if (Tnew_M > 0)
                Tnew <= Tnew_M - 1;
            else
                Tnew <= 4'h0;
        end
    end

    assign Instr_W = Instr;
    assign pc_W = pc;
    assign pc4_W = pc4;
    assign ReadData_W = ReadData;
    assign outC_W = outC;
    assign Tnew_W = Tnew;

endmodule
